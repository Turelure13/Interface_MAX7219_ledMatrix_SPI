library ieee;
use ieee.std_logic_1164.all;
library utils;
use utils.machine_state_type.all;

entity max7219 is
   
END entity;
